library verilog;
use verilog.vl_types.all;
entity Multiplex_vlg_vec_tst is
end Multiplex_vlg_vec_tst;
