library verilog;
use verilog.vl_types.all;
entity Multi21_8bits_vlg_vec_tst is
end Multi21_8bits_vlg_vec_tst;
