library verilog;
use verilog.vl_types.all;
entity HalfAdder_vlg_vec_tst is
end HalfAdder_vlg_vec_tst;
