library verilog;
use verilog.vl_types.all;
entity XOR_GATE_vlg_check_tst is
    port(
        OUTPUT          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end XOR_GATE_vlg_check_tst;
