library verilog;
use verilog.vl_types.all;
entity D_LATCH_vlg_vec_tst is
end D_LATCH_vlg_vec_tst;
