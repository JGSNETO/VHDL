library verilog;
use verilog.vl_types.all;
entity XOR_GATE_vlg_vec_tst is
end XOR_GATE_vlg_vec_tst;
