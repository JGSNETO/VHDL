library verilog;
use verilog.vl_types.all;
entity Multiplex_vlg_check_tst is
    port(
        MuxOutput       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Multiplex_vlg_check_tst;
