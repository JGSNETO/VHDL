library verilog;
use verilog.vl_types.all;
entity dff_8_vlg_vec_tst is
end dff_8_vlg_vec_tst;
