library verilog;
use verilog.vl_types.all;
entity SR_LATCH_vlg_vec_tst is
end SR_LATCH_vlg_vec_tst;
